library ieee;
  use ieee.std_logic_1164.all;
  use ieee.numeric_std.all;

entity fk is
  port (
  
  );
end entity;

architecture behavioral of fk is

begin

end architecture;
