library IEEE;
use IEEE.std_logic_1164.all;
use work.ik_pack.all;

entity cross_product is
  port (
  clock
  );
end entity;
