library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_numeric.all;

package ik_pack is
  type vec_3 is array(0 to 2) of std_logic_vector(31 downto 0);
end package;
